module CPU;
    initial $display ("Hello World.");
endmodule
