module CPU;
    initial $display (3'd6 + 3'd1);
endmodule