module CPU;
    initial $display (32'hFFFFFFF0+1);
    initial $display (32'hFFFFFFF1>>>1);
endmodule